// RTL (Verilog) generated @ Wed Mar 15 19:30:45 2017 by V3 
//               compiled @ Mar 14 2017 21:20:10
// Internal nets are renamed with prefix "v3_1489577445_".

// Module vendingMachine
module vendingMachine
(
   clk,
   reset,
   coinInNTD_50,
   coinInNTD_10,
   coinInNTD_5,
   coinInNTD_1,
   itemTypeIn,
   p,
   coinOutNTD_50,
   coinOutNTD_10,
   coinOutNTD_5,
   coinOutNTD_1,
   itemTypeOut,
   serviceTypeOut
);

   // Clock Signal for Synchronous DFF
   input clk;

   // I/O Declarations
   input reset;
   input [1:0] coinInNTD_50;
   input [1:0] coinInNTD_10;
   input [1:0] coinInNTD_5;
   input [1:0] coinInNTD_1;
   input [1:0] itemTypeIn;
   output p;
   output [2:0] coinOutNTD_50;
   output [2:0] coinOutNTD_10;
   output [2:0] coinOutNTD_5;
   output [2:0] coinOutNTD_1;
   output [1:0] itemTypeOut;
   output [1:0] serviceTypeOut;

   // Wire and Reg Declarations
   wire v3_1489577445_0;
   wire clk;
   wire reset;
   wire [1:0] coinInNTD_50;
   wire [1:0] coinInNTD_10;
   wire [1:0] coinInNTD_5;
   wire [1:0] coinInNTD_1;
   wire [1:0] itemTypeIn;
   reg [2:0] v3_1489577445_8;
   reg [2:0] v3_1489577445_9;
   reg [2:0] v3_1489577445_10;
   reg [2:0] v3_1489577445_11;
   reg [1:0] v3_1489577445_12;
   reg [1:0] v3_1489577445_13;
   reg v3_1489577445_14;
   reg [7:0] v3_1489577445_15;
   reg v3_1489577445_16;
   reg [1:0] v3_1489577445_17;
   reg [7:0] v3_1489577445_18;
   reg [2:0] v3_1489577445_19;
   reg [2:0] v3_1489577445_20;
   reg [2:0] v3_1489577445_21;
   reg [2:0] v3_1489577445_22;
   wire [2:0] v3_1489577445_23;
   wire [2:0] v3_1489577445_24;
   wire [2:0] v3_1489577445_25;
   wire [2:0] v3_1489577445_26;
   wire [2:0] v3_1489577445_27;
   wire [2:0] v3_1489577445_28;
   wire [2:0] v3_1489577445_29;
   wire [2:0] v3_1489577445_30;
   wire [2:0] v3_1489577445_31;
   wire [2:0] v3_1489577445_32;
   wire [2:0] v3_1489577445_33;
   wire [2:0] v3_1489577445_34;
   wire [2:0] v3_1489577445_35;
   wire v3_1489577445_36;
   wire v3_1489577445_37;
   wire [7:0] v3_1489577445_38;
   wire v3_1489577445_39;
   wire [1:0] v3_1489577445_40;
   wire v3_1489577445_41;
   wire [1:0] v3_1489577445_42;
   wire [2:0] v3_1489577445_43;
   wire [2:0] v3_1489577445_44;
   wire [2:0] v3_1489577445_45;
   wire [2:0] v3_1489577445_46;
   wire [2:0] v3_1489577445_47;
   wire v3_1489577445_48;
   wire v3_1489577445_49;
   wire [7:0] v3_1489577445_50;
   wire v3_1489577445_51;
   wire [1:0] v3_1489577445_52;
   wire v3_1489577445_53;
   wire [2:0] v3_1489577445_54;
   wire v3_1489577445_55;
   wire [2:0] v3_1489577445_56;
   wire [2:0] v3_1489577445_57;
   wire v3_1489577445_58;
   wire v3_1489577445_59;
   wire v3_1489577445_60;
   wire [2:0] v3_1489577445_61;
   wire v3_1489577445_62;
   wire [2:0] v3_1489577445_63;
   wire [2:0] v3_1489577445_64;
   wire [2:0] v3_1489577445_65;
   wire [2:0] v3_1489577445_66;
   wire [2:0] v3_1489577445_67;
   wire [2:0] v3_1489577445_68;
   wire [2:0] v3_1489577445_69;
   wire [2:0] v3_1489577445_70;
   wire [2:0] v3_1489577445_71;
   wire [2:0] v3_1489577445_72;
   wire [2:0] v3_1489577445_73;
   wire [2:0] v3_1489577445_74;
   wire [2:0] v3_1489577445_75;
   wire [2:0] v3_1489577445_76;
   wire [2:0] v3_1489577445_77;
   wire [2:0] v3_1489577445_78;
   wire [2:0] v3_1489577445_79;
   wire v3_1489577445_80;
   wire v3_1489577445_81;
   wire [7:0] v3_1489577445_82;
   wire [2:0] v3_1489577445_83;
   wire [2:0] v3_1489577445_84;
   wire [2:0] v3_1489577445_85;
   wire [2:0] v3_1489577445_86;
   wire [2:0] v3_1489577445_87;
   wire [2:0] v3_1489577445_88;
   wire [2:0] v3_1489577445_89;
   wire [2:0] v3_1489577445_90;
   wire [2:0] v3_1489577445_91;
   wire [2:0] v3_1489577445_92;
   wire [2:0] v3_1489577445_93;
   wire [2:0] v3_1489577445_94;
   wire [2:0] v3_1489577445_95;
   wire [2:0] v3_1489577445_96;
   wire [2:0] v3_1489577445_97;
   wire [2:0] v3_1489577445_98;
   wire [2:0] v3_1489577445_99;
   wire [2:0] v3_1489577445_100;
   wire [2:0] v3_1489577445_101;
   wire [2:0] v3_1489577445_102;
   wire [2:0] v3_1489577445_103;
   wire v3_1489577445_104;
   wire v3_1489577445_105;
   wire [7:0] v3_1489577445_106;
   wire [2:0] v3_1489577445_107;
   wire [2:0] v3_1489577445_108;
   wire [2:0] v3_1489577445_109;
   wire [2:0] v3_1489577445_110;
   wire [2:0] v3_1489577445_111;
   wire [2:0] v3_1489577445_112;
   wire [2:0] v3_1489577445_113;
   wire [2:0] v3_1489577445_114;
   wire [2:0] v3_1489577445_115;
   wire [2:0] v3_1489577445_116;
   wire [2:0] v3_1489577445_117;
   wire [2:0] v3_1489577445_118;
   wire [2:0] v3_1489577445_119;
   wire [2:0] v3_1489577445_120;
   wire [2:0] v3_1489577445_121;
   wire [2:0] v3_1489577445_122;
   wire [2:0] v3_1489577445_123;
   wire [2:0] v3_1489577445_124;
   wire [2:0] v3_1489577445_125;
   wire [2:0] v3_1489577445_126;
   wire [2:0] v3_1489577445_127;
   wire [2:0] v3_1489577445_128;
   wire [2:0] v3_1489577445_129;
   wire [2:0] v3_1489577445_130;
   wire [1:0] v3_1489577445_131;
   wire [1:0] v3_1489577445_132;
   wire [1:0] v3_1489577445_133;
   wire [1:0] v3_1489577445_134;
   wire [1:0] v3_1489577445_135;
   wire [1:0] v3_1489577445_136;
   wire [1:0] v3_1489577445_137;
   wire [1:0] v3_1489577445_138;
   wire [1:0] v3_1489577445_139;
   wire [1:0] v3_1489577445_140;
   wire [1:0] v3_1489577445_141;
   wire [1:0] v3_1489577445_142;
   wire [1:0] v3_1489577445_143;
   wire [1:0] v3_1489577445_144;
   wire v3_1489577445_145;
   wire v3_1489577445_146;
   wire [1:0] v3_1489577445_147;
   wire [1:0] v3_1489577445_148;
   wire [1:0] v3_1489577445_149;
   wire [1:0] v3_1489577445_150;
   wire [1:0] v3_1489577445_151;
   wire [1:0] v3_1489577445_152;
   wire [1:0] v3_1489577445_153;
   wire [1:0] v3_1489577445_154;
   wire [1:0] v3_1489577445_155;
   wire [1:0] v3_1489577445_156;
   wire [1:0] v3_1489577445_157;
   wire [1:0] v3_1489577445_158;
   wire [1:0] v3_1489577445_159;
   wire [1:0] v3_1489577445_160;
   wire [1:0] v3_1489577445_161;
   wire [1:0] v3_1489577445_162;
   wire [1:0] v3_1489577445_163;
   wire [1:0] v3_1489577445_164;
   wire [1:0] v3_1489577445_165;
   wire [1:0] v3_1489577445_166;
   wire [1:0] v3_1489577445_167;
   wire [1:0] v3_1489577445_168;
   wire [1:0] v3_1489577445_169;
   wire v3_1489577445_170;
   wire v3_1489577445_171;
   wire v3_1489577445_172;
   wire v3_1489577445_173;
   wire v3_1489577445_174;
   wire [7:0] v3_1489577445_175;
   wire [7:0] v3_1489577445_176;
   wire [7:0] v3_1489577445_177;
   wire [7:0] v3_1489577445_178;
   wire [7:0] v3_1489577445_179;
   wire [7:0] v3_1489577445_180;
   wire [7:0] v3_1489577445_181;
   wire [7:0] v3_1489577445_182;
   wire [7:0] v3_1489577445_183;
   wire [7:0] v3_1489577445_184;
   wire [5:0] v3_1489577445_185;
   wire [7:0] v3_1489577445_186;
   wire [7:0] v3_1489577445_187;
   wire [7:0] v3_1489577445_188;
   wire [7:0] v3_1489577445_189;
   wire [7:0] v3_1489577445_190;
   wire [7:0] v3_1489577445_191;
   wire [7:0] v3_1489577445_192;
   wire [7:0] v3_1489577445_193;
   wire [7:0] v3_1489577445_194;
   wire [7:0] v3_1489577445_195;
   wire [7:0] v3_1489577445_196;
   wire [7:0] v3_1489577445_197;
   wire [7:0] v3_1489577445_198;
   wire [7:0] v3_1489577445_199;
   wire [7:0] v3_1489577445_200;
   wire [7:0] v3_1489577445_201;
   wire [7:0] v3_1489577445_202;
   wire [7:0] v3_1489577445_203;
   wire [7:0] v3_1489577445_204;
   wire [7:0] v3_1489577445_205;
   wire v3_1489577445_206;
   wire v3_1489577445_207;
   wire v3_1489577445_208;
   wire v3_1489577445_209;
   wire v3_1489577445_210;
   wire v3_1489577445_211;
   wire v3_1489577445_212;
   wire v3_1489577445_213;
   wire v3_1489577445_214;
   wire v3_1489577445_215;
   wire v3_1489577445_216;
   wire v3_1489577445_217;
   wire v3_1489577445_218;
   wire v3_1489577445_219;
   wire [1:0] v3_1489577445_220;
   wire [1:0] v3_1489577445_221;
   wire [1:0] v3_1489577445_222;
   wire [1:0] v3_1489577445_223;
   wire [1:0] v3_1489577445_224;
   wire [1:0] v3_1489577445_225;
   wire [1:0] v3_1489577445_226;
   wire [1:0] v3_1489577445_227;
   wire [1:0] v3_1489577445_228;
   wire [1:0] v3_1489577445_229;
   wire [1:0] v3_1489577445_230;
   wire [1:0] v3_1489577445_231;
   wire [1:0] v3_1489577445_232;
   wire [1:0] v3_1489577445_233;
   wire [1:0] v3_1489577445_234;
   wire [1:0] v3_1489577445_235;
   wire [1:0] v3_1489577445_236;
   wire [1:0] v3_1489577445_237;
   wire [1:0] v3_1489577445_238;
   wire [1:0] v3_1489577445_239;
   wire [1:0] v3_1489577445_240;
   wire [1:0] v3_1489577445_241;
   wire [1:0] v3_1489577445_242;
   wire [1:0] v3_1489577445_243;
   wire [1:0] v3_1489577445_244;
   wire [1:0] v3_1489577445_245;
   wire [1:0] v3_1489577445_246;
   wire [1:0] v3_1489577445_247;
   wire [1:0] v3_1489577445_248;
   wire [7:0] v3_1489577445_249;
   wire [7:0] v3_1489577445_250;
   wire [7:0] v3_1489577445_251;
   wire [7:0] v3_1489577445_252;
   wire [7:0] v3_1489577445_253;
   wire [7:0] v3_1489577445_254;
   wire [7:0] v3_1489577445_255;
   wire [7:0] v3_1489577445_256;
   wire [7:0] v3_1489577445_257;
   wire [7:0] v3_1489577445_258;
   wire [7:0] v3_1489577445_259;
   wire [7:0] v3_1489577445_260;
   wire [7:0] v3_1489577445_261;
   wire [7:0] v3_1489577445_262;
   wire [7:0] v3_1489577445_263;
   wire [7:0] v3_1489577445_264;
   wire [7:0] v3_1489577445_265;
   wire [7:0] v3_1489577445_266;
   wire [7:0] v3_1489577445_267;
   wire [7:0] v3_1489577445_268;
   wire [7:0] v3_1489577445_269;
   wire [7:0] v3_1489577445_270;
   wire [7:0] v3_1489577445_271;
   wire [7:0] v3_1489577445_272;
   wire [7:0] v3_1489577445_273;
   wire [7:0] v3_1489577445_274;
   wire [7:0] v3_1489577445_275;
   wire [7:0] v3_1489577445_276;
   wire [7:0] v3_1489577445_277;
   wire [7:0] v3_1489577445_278;
   wire [7:0] v3_1489577445_279;
   wire [7:0] v3_1489577445_280;
   wire [7:0] v3_1489577445_281;
   wire [7:0] v3_1489577445_282;
   wire [7:0] v3_1489577445_283;
   wire v3_1489577445_284;
   wire [7:0] v3_1489577445_285;
   wire v3_1489577445_286;
   wire [7:0] v3_1489577445_287;
   wire v3_1489577445_288;
   wire [7:0] v3_1489577445_289;
   wire [7:0] v3_1489577445_290;
   wire [2:0] v3_1489577445_291;
   wire [2:0] v3_1489577445_292;
   wire [2:0] v3_1489577445_293;
   wire [2:0] v3_1489577445_294;
   wire [2:0] v3_1489577445_295;
   wire [2:0] v3_1489577445_296;
   wire [2:0] v3_1489577445_297;
   wire [2:0] v3_1489577445_298;
   wire [2:0] v3_1489577445_299;
   wire [2:0] v3_1489577445_300;
   wire [2:0] v3_1489577445_301;
   wire [2:0] v3_1489577445_302;
   wire [2:0] v3_1489577445_303;
   wire [2:0] v3_1489577445_304;
   wire [2:0] v3_1489577445_305;
   wire [2:0] v3_1489577445_306;
   wire [2:0] v3_1489577445_307;
   wire [2:0] v3_1489577445_308;
   wire [2:0] v3_1489577445_309;
   wire [2:0] v3_1489577445_310;
   wire [2:0] v3_1489577445_311;
   wire [2:0] v3_1489577445_312;
   wire [2:0] v3_1489577445_313;
   wire [2:0] v3_1489577445_314;
   wire v3_1489577445_315;
   wire [3:0] v3_1489577445_316;
   wire [3:0] v3_1489577445_317;
   wire [3:0] v3_1489577445_318;
   wire [3:0] v3_1489577445_319;
   wire [3:0] v3_1489577445_320;
   wire [3:0] v3_1489577445_321;
   wire [3:0] v3_1489577445_322;
   wire [2:0] v3_1489577445_323;
   wire [2:0] v3_1489577445_324;
   wire [2:0] v3_1489577445_325;
   wire [2:0] v3_1489577445_326;
   wire [2:0] v3_1489577445_327;
   wire [2:0] v3_1489577445_328;
   wire [2:0] v3_1489577445_329;
   wire [2:0] v3_1489577445_330;
   wire [2:0] v3_1489577445_331;
   wire [2:0] v3_1489577445_332;
   wire [2:0] v3_1489577445_333;
   wire [2:0] v3_1489577445_334;
   wire [2:0] v3_1489577445_335;
   wire [2:0] v3_1489577445_336;
   wire [2:0] v3_1489577445_337;
   wire [2:0] v3_1489577445_338;
   wire [2:0] v3_1489577445_339;
   wire [2:0] v3_1489577445_340;
   wire [2:0] v3_1489577445_341;
   wire [2:0] v3_1489577445_342;
   wire [2:0] v3_1489577445_343;
   wire [2:0] v3_1489577445_344;
   wire [2:0] v3_1489577445_345;
   wire [2:0] v3_1489577445_346;
   wire [2:0] v3_1489577445_347;
   wire [2:0] v3_1489577445_348;
   wire v3_1489577445_349;
   wire [3:0] v3_1489577445_350;
   wire [3:0] v3_1489577445_351;
   wire [3:0] v3_1489577445_352;
   wire [3:0] v3_1489577445_353;
   wire [3:0] v3_1489577445_354;
   wire [3:0] v3_1489577445_355;
   wire [2:0] v3_1489577445_356;
   wire [2:0] v3_1489577445_357;
   wire [2:0] v3_1489577445_358;
   wire [2:0] v3_1489577445_359;
   wire [2:0] v3_1489577445_360;
   wire [2:0] v3_1489577445_361;
   wire [2:0] v3_1489577445_362;
   wire [2:0] v3_1489577445_363;
   wire [2:0] v3_1489577445_364;
   wire [2:0] v3_1489577445_365;
   wire [2:0] v3_1489577445_366;
   wire [2:0] v3_1489577445_367;
   wire [2:0] v3_1489577445_368;
   wire [2:0] v3_1489577445_369;
   wire [2:0] v3_1489577445_370;
   wire [2:0] v3_1489577445_371;
   wire [2:0] v3_1489577445_372;
   wire [2:0] v3_1489577445_373;
   wire [2:0] v3_1489577445_374;
   wire [2:0] v3_1489577445_375;
   wire [2:0] v3_1489577445_376;
   wire [2:0] v3_1489577445_377;
   wire [2:0] v3_1489577445_378;
   wire v3_1489577445_379;
   wire [3:0] v3_1489577445_380;
   wire [3:0] v3_1489577445_381;
   wire [3:0] v3_1489577445_382;
   wire [3:0] v3_1489577445_383;
   wire [3:0] v3_1489577445_384;
   wire [3:0] v3_1489577445_385;
   wire [2:0] v3_1489577445_386;
   wire [2:0] v3_1489577445_387;
   wire [2:0] v3_1489577445_388;
   wire [2:0] v3_1489577445_389;
   wire [2:0] v3_1489577445_390;
   wire [2:0] v3_1489577445_391;
   wire [2:0] v3_1489577445_392;
   wire [2:0] v3_1489577445_393;
   wire [2:0] v3_1489577445_394;
   wire [2:0] v3_1489577445_395;
   wire [2:0] v3_1489577445_396;
   wire [2:0] v3_1489577445_397;
   wire [2:0] v3_1489577445_398;
   wire [2:0] v3_1489577445_399;
   wire [2:0] v3_1489577445_400;
   wire [2:0] v3_1489577445_401;
   wire [2:0] v3_1489577445_402;
   wire [2:0] v3_1489577445_403;
   wire [2:0] v3_1489577445_404;
   wire [2:0] v3_1489577445_405;
   wire [2:0] v3_1489577445_406;
   wire [2:0] v3_1489577445_407;
   wire [2:0] v3_1489577445_408;
   wire [2:0] v3_1489577445_409;
   wire [2:0] v3_1489577445_410;
   wire v3_1489577445_411;
   wire [3:0] v3_1489577445_412;
   wire [3:0] v3_1489577445_413;
   wire [3:0] v3_1489577445_414;
   wire [3:0] v3_1489577445_415;
   wire [3:0] v3_1489577445_416;
   wire [3:0] v3_1489577445_417;
   wire [2:0] v3_1489577445_418;
   wire [2:0] v3_1489577445_419;
   wire v3_1489577445_420;
   wire v3_1489577445_421;
   wire v3_1489577445_422;
   wire v3_1489577445_423;
   wire v3_1489577445_424;
   wire v3_1489577445_425;
   wire v3_1489577445_426;
   wire v3_1489577445_427;
   wire [7:0] v3_1489577445_428;
   wire [7:0] v3_1489577445_429;
   wire [7:0] v3_1489577445_430;
   wire [7:0] v3_1489577445_431;
   wire [7:0] v3_1489577445_432;
   wire [4:0] v3_1489577445_433;
   wire [7:0] v3_1489577445_434;
   wire [7:0] v3_1489577445_435;
   wire [7:0] v3_1489577445_436;
   wire [7:0] v3_1489577445_437;
   wire [7:0] v3_1489577445_438;
   wire [7:0] v3_1489577445_439;
   wire [7:0] v3_1489577445_440;
   wire [7:0] v3_1489577445_441;
   wire [7:0] v3_1489577445_442;
   wire [7:0] v3_1489577445_443;
   wire [7:0] v3_1489577445_444;
   wire [7:0] v3_1489577445_445;
   wire [7:0] v3_1489577445_446;
   wire [7:0] v3_1489577445_447;
   wire [7:0] v3_1489577445_448;
   wire [7:0] v3_1489577445_449;
   wire [7:0] v3_1489577445_450;
   wire v3_1489577445_451;

   // Output Net Declarations
   wire p;
   wire [2:0] coinOutNTD_50;
   wire [2:0] coinOutNTD_10;
   wire [2:0] coinOutNTD_5;
   wire [2:0] coinOutNTD_1;
   wire [1:0] itemTypeOut;
   wire [1:0] serviceTypeOut;

   // Combinational Assignments
   assign v3_1489577445_0 = 1'b0; 
   assign v3_1489577445_23 = v3_1489577445_62 ? v3_1489577445_61 : v3_1489577445_24;
   assign v3_1489577445_24 = v3_1489577445_25;
   assign v3_1489577445_25 = v3_1489577445_60 ? v3_1489577445_56 : v3_1489577445_26;
   assign v3_1489577445_26 = v3_1489577445_55 ? v3_1489577445_54 : v3_1489577445_27;
   assign v3_1489577445_27 = v3_1489577445_53 ? v3_1489577445_32 : v3_1489577445_28;
   assign v3_1489577445_28 = v3_1489577445_51 ? v3_1489577445_43 : v3_1489577445_29;
   assign v3_1489577445_29 = v3_1489577445_41 ? v3_1489577445_32 : v3_1489577445_30;
   assign v3_1489577445_30 = v3_1489577445_39 ? v3_1489577445_32 : v3_1489577445_31;
   assign v3_1489577445_31 = v3_1489577445_37 ? v3_1489577445_33 : v3_1489577445_32;
   assign v3_1489577445_32 = v3_1489577445_8;
   assign v3_1489577445_33 = v3_1489577445_36 ? v3_1489577445_34 : v3_1489577445_32;
   assign v3_1489577445_34 = v3_1489577445_35;
   assign v3_1489577445_35 = 3'b000; 
   assign v3_1489577445_36 = v3_1489577445_21 == v3_1489577445_35;
   assign v3_1489577445_37 = v3_1489577445_18 >= v3_1489577445_38;
   assign v3_1489577445_38 = 8'b00000001; 
   assign v3_1489577445_39 = v3_1489577445_17 == v3_1489577445_40;
   assign v3_1489577445_40 = 2'b10; 
   assign v3_1489577445_41 = v3_1489577445_17 == v3_1489577445_42;
   assign v3_1489577445_42 = 2'b01; 
   assign v3_1489577445_43 = v3_1489577445_49 ? v3_1489577445_44 : v3_1489577445_32;
   assign v3_1489577445_44 = v3_1489577445_48 ? v3_1489577445_32 : v3_1489577445_45;
   assign v3_1489577445_45 = v3_1489577445_47;
   assign v3_1489577445_46 = 3'b001; 
   assign v3_1489577445_47 = v3_1489577445_8 + v3_1489577445_46;
   assign v3_1489577445_48 = v3_1489577445_19 == v3_1489577445_35;
   assign v3_1489577445_49 = v3_1489577445_18 >= v3_1489577445_50;
   assign v3_1489577445_50 = 8'b00110010; 
   assign v3_1489577445_51 = v3_1489577445_17 == v3_1489577445_52;
   assign v3_1489577445_52 = 2'b00; 
   assign v3_1489577445_53 = ~v3_1489577445_16;
   assign v3_1489577445_54 = v3_1489577445_35;
   assign v3_1489577445_55 = v3_1489577445_13 == v3_1489577445_52;
   assign v3_1489577445_56 = v3_1489577445_58 ? v3_1489577445_57 : v3_1489577445_32;
   assign v3_1489577445_57 = v3_1489577445_35;
   assign v3_1489577445_58 = ~v3_1489577445_59;
   assign v3_1489577445_59 = itemTypeIn == v3_1489577445_52;
   assign v3_1489577445_60 = v3_1489577445_13 == v3_1489577445_42;
   assign v3_1489577445_61 = v3_1489577445_35;
   assign v3_1489577445_62 = ~reset;
   assign v3_1489577445_63 = 3'b000; 
   assign v3_1489577445_64 = v3_1489577445_62 ? v3_1489577445_86 : v3_1489577445_65;
   assign v3_1489577445_65 = v3_1489577445_66;
   assign v3_1489577445_66 = v3_1489577445_60 ? v3_1489577445_84 : v3_1489577445_67;
   assign v3_1489577445_67 = v3_1489577445_55 ? v3_1489577445_83 : v3_1489577445_68;
   assign v3_1489577445_68 = v3_1489577445_53 ? v3_1489577445_73 : v3_1489577445_69;
   assign v3_1489577445_69 = v3_1489577445_51 ? v3_1489577445_73 : v3_1489577445_70;
   assign v3_1489577445_70 = v3_1489577445_41 ? v3_1489577445_76 : v3_1489577445_71;
   assign v3_1489577445_71 = v3_1489577445_39 ? v3_1489577445_73 : v3_1489577445_72;
   assign v3_1489577445_72 = v3_1489577445_37 ? v3_1489577445_74 : v3_1489577445_73;
   assign v3_1489577445_73 = v3_1489577445_9;
   assign v3_1489577445_74 = v3_1489577445_36 ? v3_1489577445_75 : v3_1489577445_73;
   assign v3_1489577445_75 = v3_1489577445_35;
   assign v3_1489577445_76 = v3_1489577445_81 ? v3_1489577445_77 : v3_1489577445_73;
   assign v3_1489577445_77 = v3_1489577445_80 ? v3_1489577445_73 : v3_1489577445_78;
   assign v3_1489577445_78 = v3_1489577445_79;
   assign v3_1489577445_79 = v3_1489577445_9 + v3_1489577445_46;
   assign v3_1489577445_80 = v3_1489577445_20 == v3_1489577445_35;
   assign v3_1489577445_81 = v3_1489577445_18 >= v3_1489577445_82;
   assign v3_1489577445_82 = 8'b00001010; 
   assign v3_1489577445_83 = v3_1489577445_35;
   assign v3_1489577445_84 = v3_1489577445_58 ? v3_1489577445_85 : v3_1489577445_73;
   assign v3_1489577445_85 = v3_1489577445_35;
   assign v3_1489577445_86 = v3_1489577445_35;
   assign v3_1489577445_87 = 3'b000; 
   assign v3_1489577445_88 = v3_1489577445_62 ? v3_1489577445_110 : v3_1489577445_89;
   assign v3_1489577445_89 = v3_1489577445_90;
   assign v3_1489577445_90 = v3_1489577445_60 ? v3_1489577445_108 : v3_1489577445_91;
   assign v3_1489577445_91 = v3_1489577445_55 ? v3_1489577445_107 : v3_1489577445_92;
   assign v3_1489577445_92 = v3_1489577445_53 ? v3_1489577445_97 : v3_1489577445_93;
   assign v3_1489577445_93 = v3_1489577445_51 ? v3_1489577445_97 : v3_1489577445_94;
   assign v3_1489577445_94 = v3_1489577445_41 ? v3_1489577445_97 : v3_1489577445_95;
   assign v3_1489577445_95 = v3_1489577445_39 ? v3_1489577445_100 : v3_1489577445_96;
   assign v3_1489577445_96 = v3_1489577445_37 ? v3_1489577445_98 : v3_1489577445_97;
   assign v3_1489577445_97 = v3_1489577445_10;
   assign v3_1489577445_98 = v3_1489577445_36 ? v3_1489577445_99 : v3_1489577445_97;
   assign v3_1489577445_99 = v3_1489577445_35;
   assign v3_1489577445_100 = v3_1489577445_105 ? v3_1489577445_101 : v3_1489577445_97;
   assign v3_1489577445_101 = v3_1489577445_104 ? v3_1489577445_97 : v3_1489577445_102;
   assign v3_1489577445_102 = v3_1489577445_103;
   assign v3_1489577445_103 = v3_1489577445_10 + v3_1489577445_46;
   assign v3_1489577445_104 = v3_1489577445_22 == v3_1489577445_35;
   assign v3_1489577445_105 = v3_1489577445_18 >= v3_1489577445_106;
   assign v3_1489577445_106 = 8'b00000101; 
   assign v3_1489577445_107 = v3_1489577445_35;
   assign v3_1489577445_108 = v3_1489577445_58 ? v3_1489577445_109 : v3_1489577445_97;
   assign v3_1489577445_109 = v3_1489577445_35;
   assign v3_1489577445_110 = v3_1489577445_35;
   assign v3_1489577445_111 = 3'b000; 
   assign v3_1489577445_112 = v3_1489577445_62 ? v3_1489577445_129 : v3_1489577445_113;
   assign v3_1489577445_113 = v3_1489577445_114;
   assign v3_1489577445_114 = v3_1489577445_60 ? v3_1489577445_127 : v3_1489577445_115;
   assign v3_1489577445_115 = v3_1489577445_55 ? v3_1489577445_126 : v3_1489577445_116;
   assign v3_1489577445_116 = v3_1489577445_53 ? v3_1489577445_121 : v3_1489577445_117;
   assign v3_1489577445_117 = v3_1489577445_51 ? v3_1489577445_121 : v3_1489577445_118;
   assign v3_1489577445_118 = v3_1489577445_41 ? v3_1489577445_121 : v3_1489577445_119;
   assign v3_1489577445_119 = v3_1489577445_39 ? v3_1489577445_121 : v3_1489577445_120;
   assign v3_1489577445_120 = v3_1489577445_37 ? v3_1489577445_122 : v3_1489577445_121;
   assign v3_1489577445_121 = v3_1489577445_11;
   assign v3_1489577445_122 = v3_1489577445_36 ? v3_1489577445_125 : v3_1489577445_123;
   assign v3_1489577445_123 = v3_1489577445_124;
   assign v3_1489577445_124 = v3_1489577445_11 + v3_1489577445_46;
   assign v3_1489577445_125 = v3_1489577445_35;
   assign v3_1489577445_126 = v3_1489577445_35;
   assign v3_1489577445_127 = v3_1489577445_58 ? v3_1489577445_128 : v3_1489577445_121;
   assign v3_1489577445_128 = v3_1489577445_35;
   assign v3_1489577445_129 = v3_1489577445_35;
   assign v3_1489577445_130 = 3'b000; 
   assign v3_1489577445_131 = v3_1489577445_62 ? v3_1489577445_150 : v3_1489577445_132;
   assign v3_1489577445_132 = v3_1489577445_133;
   assign v3_1489577445_133 = v3_1489577445_60 ? v3_1489577445_148 : v3_1489577445_134;
   assign v3_1489577445_134 = v3_1489577445_55 ? v3_1489577445_147 : v3_1489577445_135;
   assign v3_1489577445_135 = v3_1489577445_53 ? v3_1489577445_143 : v3_1489577445_136;
   assign v3_1489577445_136 = v3_1489577445_51 ? v3_1489577445_140 : v3_1489577445_137;
   assign v3_1489577445_137 = v3_1489577445_41 ? v3_1489577445_140 : v3_1489577445_138;
   assign v3_1489577445_138 = v3_1489577445_39 ? v3_1489577445_140 : v3_1489577445_139;
   assign v3_1489577445_139 = v3_1489577445_37 ? v3_1489577445_141 : v3_1489577445_140;
   assign v3_1489577445_140 = v3_1489577445_12;
   assign v3_1489577445_141 = v3_1489577445_36 ? v3_1489577445_142 : v3_1489577445_140;
   assign v3_1489577445_142 = v3_1489577445_52;
   assign v3_1489577445_143 = v3_1489577445_145 ? v3_1489577445_144 : v3_1489577445_140;
   assign v3_1489577445_144 = v3_1489577445_52;
   assign v3_1489577445_145 = ~v3_1489577445_146;
   assign v3_1489577445_146 = v3_1489577445_15 >= v3_1489577445_18;
   assign v3_1489577445_147 = v3_1489577445_52;
   assign v3_1489577445_148 = v3_1489577445_58 ? v3_1489577445_149 : v3_1489577445_140;
   assign v3_1489577445_149 = itemTypeIn;
   assign v3_1489577445_150 = v3_1489577445_52;
   assign v3_1489577445_151 = 2'b00; 
   assign v3_1489577445_152 = v3_1489577445_62 ? v3_1489577445_168 : v3_1489577445_153;
   assign v3_1489577445_153 = v3_1489577445_154;
   assign v3_1489577445_154 = v3_1489577445_60 ? v3_1489577445_166 : v3_1489577445_155;
   assign v3_1489577445_155 = v3_1489577445_55 ? v3_1489577445_165 : v3_1489577445_156;
   assign v3_1489577445_156 = v3_1489577445_53 ? v3_1489577445_163 : v3_1489577445_157;
   assign v3_1489577445_157 = v3_1489577445_51 ? v3_1489577445_163 : v3_1489577445_158;
   assign v3_1489577445_158 = v3_1489577445_41 ? v3_1489577445_163 : v3_1489577445_159;
   assign v3_1489577445_159 = v3_1489577445_39 ? v3_1489577445_163 : v3_1489577445_160;
   assign v3_1489577445_160 = v3_1489577445_37 ? v3_1489577445_162 : v3_1489577445_161;
   assign v3_1489577445_161 = v3_1489577445_52;
   assign v3_1489577445_162 = v3_1489577445_36 ? v3_1489577445_164 : v3_1489577445_163;
   assign v3_1489577445_163 = v3_1489577445_13;
   assign v3_1489577445_164 = v3_1489577445_52;
   assign v3_1489577445_165 = v3_1489577445_42;
   assign v3_1489577445_166 = v3_1489577445_58 ? v3_1489577445_167 : v3_1489577445_163;
   assign v3_1489577445_167 = v3_1489577445_40;
   assign v3_1489577445_168 = v3_1489577445_42;
   assign v3_1489577445_169 = 2'b00; 
   assign v3_1489577445_170 = v3_1489577445_62 ? v3_1489577445_172 : v3_1489577445_171;
   assign v3_1489577445_171 = v3_1489577445_14;
   assign v3_1489577445_172 = v3_1489577445_173;
   assign v3_1489577445_173 = 1'b1; 
   assign v3_1489577445_174 = 1'b0; 
   assign v3_1489577445_175 = v3_1489577445_62 ? v3_1489577445_203 : v3_1489577445_176;
   assign v3_1489577445_176 = v3_1489577445_177;
   assign v3_1489577445_177 = v3_1489577445_60 ? v3_1489577445_179 : v3_1489577445_178;
   assign v3_1489577445_178 = v3_1489577445_15;
   assign v3_1489577445_179 = v3_1489577445_58 ? v3_1489577445_180 : v3_1489577445_178;
   assign v3_1489577445_180 = v3_1489577445_202;
   assign v3_1489577445_181 = v3_1489577445_197;
   assign v3_1489577445_182 = v3_1489577445_192;
   assign v3_1489577445_183 = v3_1489577445_187;
   assign v3_1489577445_184 = v3_1489577445_186;
   assign v3_1489577445_185 = 6'b000000; 
   assign v3_1489577445_186 = {v3_1489577445_185, coinInNTD_50};
   assign v3_1489577445_187 = v3_1489577445_50 * v3_1489577445_184;
   assign v3_1489577445_188 = v3_1489577445_191;
   assign v3_1489577445_189 = v3_1489577445_190;
   assign v3_1489577445_190 = {v3_1489577445_185, coinInNTD_10};
   assign v3_1489577445_191 = v3_1489577445_82 * v3_1489577445_189;
   assign v3_1489577445_192 = v3_1489577445_183 + v3_1489577445_188;
   assign v3_1489577445_193 = v3_1489577445_196;
   assign v3_1489577445_194 = v3_1489577445_195;
   assign v3_1489577445_195 = {v3_1489577445_185, coinInNTD_5};
   assign v3_1489577445_196 = v3_1489577445_106 * v3_1489577445_194;
   assign v3_1489577445_197 = v3_1489577445_182 + v3_1489577445_193;
   assign v3_1489577445_198 = v3_1489577445_201;
   assign v3_1489577445_199 = v3_1489577445_200;
   assign v3_1489577445_200 = {v3_1489577445_185, coinInNTD_1};
   assign v3_1489577445_201 = v3_1489577445_38 * v3_1489577445_199;
   assign v3_1489577445_202 = v3_1489577445_181 + v3_1489577445_198;
   assign v3_1489577445_203 = v3_1489577445_204;
   assign v3_1489577445_204 = 8'b00000000; 
   assign v3_1489577445_205 = 8'b00000000; 
   assign v3_1489577445_206 = v3_1489577445_62 ? v3_1489577445_218 : v3_1489577445_207;
   assign v3_1489577445_207 = v3_1489577445_208;
   assign v3_1489577445_208 = v3_1489577445_60 ? v3_1489577445_215 : v3_1489577445_209;
   assign v3_1489577445_209 = v3_1489577445_55 ? v3_1489577445_211 : v3_1489577445_210;
   assign v3_1489577445_210 = v3_1489577445_53 ? v3_1489577445_212 : v3_1489577445_211;
   assign v3_1489577445_211 = v3_1489577445_16;
   assign v3_1489577445_212 = v3_1489577445_145 ? v3_1489577445_214 : v3_1489577445_213;
   assign v3_1489577445_213 = v3_1489577445_173;
   assign v3_1489577445_214 = v3_1489577445_173;
   assign v3_1489577445_215 = v3_1489577445_58 ? v3_1489577445_216 : v3_1489577445_211;
   assign v3_1489577445_216 = v3_1489577445_217;
   assign v3_1489577445_217 = 1'b0; 
   assign v3_1489577445_218 = v3_1489577445_217;
   assign v3_1489577445_219 = 1'b0; 
   assign v3_1489577445_220 = v3_1489577445_62 ? v3_1489577445_247 : v3_1489577445_221;
   assign v3_1489577445_221 = v3_1489577445_222;
   assign v3_1489577445_222 = v3_1489577445_60 ? v3_1489577445_245 : v3_1489577445_223;
   assign v3_1489577445_223 = v3_1489577445_55 ? v3_1489577445_229 : v3_1489577445_224;
   assign v3_1489577445_224 = v3_1489577445_53 ? v3_1489577445_229 : v3_1489577445_225;
   assign v3_1489577445_225 = v3_1489577445_51 ? v3_1489577445_241 : v3_1489577445_226;
   assign v3_1489577445_226 = v3_1489577445_41 ? v3_1489577445_237 : v3_1489577445_227;
   assign v3_1489577445_227 = v3_1489577445_39 ? v3_1489577445_232 : v3_1489577445_228;
   assign v3_1489577445_228 = v3_1489577445_37 ? v3_1489577445_230 : v3_1489577445_229;
   assign v3_1489577445_229 = v3_1489577445_17;
   assign v3_1489577445_230 = v3_1489577445_36 ? v3_1489577445_231 : v3_1489577445_229;
   assign v3_1489577445_231 = v3_1489577445_52;
   assign v3_1489577445_232 = v3_1489577445_105 ? v3_1489577445_235 : v3_1489577445_233;
   assign v3_1489577445_233 = v3_1489577445_234;
   assign v3_1489577445_234 = 2'b11; 
   assign v3_1489577445_235 = v3_1489577445_104 ? v3_1489577445_236 : v3_1489577445_229;
   assign v3_1489577445_236 = v3_1489577445_234;
   assign v3_1489577445_237 = v3_1489577445_81 ? v3_1489577445_239 : v3_1489577445_238;
   assign v3_1489577445_238 = v3_1489577445_40;
   assign v3_1489577445_239 = v3_1489577445_80 ? v3_1489577445_240 : v3_1489577445_229;
   assign v3_1489577445_240 = v3_1489577445_40;
   assign v3_1489577445_241 = v3_1489577445_49 ? v3_1489577445_243 : v3_1489577445_242;
   assign v3_1489577445_242 = v3_1489577445_42;
   assign v3_1489577445_243 = v3_1489577445_48 ? v3_1489577445_244 : v3_1489577445_229;
   assign v3_1489577445_244 = v3_1489577445_42;
   assign v3_1489577445_245 = v3_1489577445_58 ? v3_1489577445_246 : v3_1489577445_229;
   assign v3_1489577445_246 = v3_1489577445_52;
   assign v3_1489577445_247 = v3_1489577445_52;
   assign v3_1489577445_248 = 2'b00; 
   assign v3_1489577445_249 = v3_1489577445_62 ? v3_1489577445_289 : v3_1489577445_250;
   assign v3_1489577445_250 = v3_1489577445_251;
   assign v3_1489577445_251 = v3_1489577445_60 ? v3_1489577445_279 : v3_1489577445_252;
   assign v3_1489577445_252 = v3_1489577445_55 ? v3_1489577445_258 : v3_1489577445_253;
   assign v3_1489577445_253 = v3_1489577445_53 ? v3_1489577445_275 : v3_1489577445_254;
   assign v3_1489577445_254 = v3_1489577445_51 ? v3_1489577445_271 : v3_1489577445_255;
   assign v3_1489577445_255 = v3_1489577445_41 ? v3_1489577445_267 : v3_1489577445_256;
   assign v3_1489577445_256 = v3_1489577445_39 ? v3_1489577445_263 : v3_1489577445_257;
   assign v3_1489577445_257 = v3_1489577445_37 ? v3_1489577445_259 : v3_1489577445_258;
   assign v3_1489577445_258 = v3_1489577445_18;
   assign v3_1489577445_259 = v3_1489577445_36 ? v3_1489577445_262 : v3_1489577445_260;
   assign v3_1489577445_260 = v3_1489577445_261;
   assign v3_1489577445_261 = v3_1489577445_18 - v3_1489577445_38;
   assign v3_1489577445_262 = v3_1489577445_15;
   assign v3_1489577445_263 = v3_1489577445_105 ? v3_1489577445_264 : v3_1489577445_258;
   assign v3_1489577445_264 = v3_1489577445_104 ? v3_1489577445_258 : v3_1489577445_265;
   assign v3_1489577445_265 = v3_1489577445_266;
   assign v3_1489577445_266 = v3_1489577445_18 - v3_1489577445_106;
   assign v3_1489577445_267 = v3_1489577445_81 ? v3_1489577445_268 : v3_1489577445_258;
   assign v3_1489577445_268 = v3_1489577445_80 ? v3_1489577445_258 : v3_1489577445_269;
   assign v3_1489577445_269 = v3_1489577445_270;
   assign v3_1489577445_270 = v3_1489577445_18 - v3_1489577445_82;
   assign v3_1489577445_271 = v3_1489577445_49 ? v3_1489577445_272 : v3_1489577445_258;
   assign v3_1489577445_272 = v3_1489577445_48 ? v3_1489577445_258 : v3_1489577445_273;
   assign v3_1489577445_273 = v3_1489577445_274;
   assign v3_1489577445_274 = v3_1489577445_18 - v3_1489577445_50;
   assign v3_1489577445_275 = v3_1489577445_145 ? v3_1489577445_278 : v3_1489577445_276;
   assign v3_1489577445_276 = v3_1489577445_277;
   assign v3_1489577445_277 = v3_1489577445_15 - v3_1489577445_18;
   assign v3_1489577445_278 = v3_1489577445_15;
   assign v3_1489577445_279 = v3_1489577445_58 ? v3_1489577445_280 : v3_1489577445_258;
   assign v3_1489577445_280 = v3_1489577445_288 ? v3_1489577445_287 : v3_1489577445_281;
   assign v3_1489577445_281 = v3_1489577445_286 ? v3_1489577445_285 : v3_1489577445_282;
   assign v3_1489577445_282 = v3_1489577445_284 ? v3_1489577445_283 : v3_1489577445_204;
   assign v3_1489577445_283 = 8'b00010110; 
   assign v3_1489577445_284 = itemTypeIn == v3_1489577445_234;
   assign v3_1489577445_285 = 8'b00001111; 
   assign v3_1489577445_286 = itemTypeIn == v3_1489577445_40;
   assign v3_1489577445_287 = 8'b00001000; 
   assign v3_1489577445_288 = itemTypeIn == v3_1489577445_42;
   assign v3_1489577445_289 = v3_1489577445_204;
   assign v3_1489577445_290 = 8'b00000000; 
   assign v3_1489577445_291 = v3_1489577445_62 ? v3_1489577445_323 : v3_1489577445_292;
   assign v3_1489577445_292 = v3_1489577445_293;
   assign v3_1489577445_293 = v3_1489577445_60 ? v3_1489577445_308 : v3_1489577445_294;
   assign v3_1489577445_294 = v3_1489577445_55 ? v3_1489577445_300 : v3_1489577445_295;
   assign v3_1489577445_295 = v3_1489577445_53 ? v3_1489577445_300 : v3_1489577445_296;
   assign v3_1489577445_296 = v3_1489577445_51 ? v3_1489577445_304 : v3_1489577445_297;
   assign v3_1489577445_297 = v3_1489577445_41 ? v3_1489577445_300 : v3_1489577445_298;
   assign v3_1489577445_298 = v3_1489577445_39 ? v3_1489577445_300 : v3_1489577445_299;
   assign v3_1489577445_299 = v3_1489577445_37 ? v3_1489577445_301 : v3_1489577445_300;
   assign v3_1489577445_300 = v3_1489577445_19;
   assign v3_1489577445_301 = v3_1489577445_36 ? v3_1489577445_302 : v3_1489577445_300;
   assign v3_1489577445_302 = v3_1489577445_303;
   assign v3_1489577445_303 = v3_1489577445_19 + v3_1489577445_8;
   assign v3_1489577445_304 = v3_1489577445_49 ? v3_1489577445_305 : v3_1489577445_300;
   assign v3_1489577445_305 = v3_1489577445_48 ? v3_1489577445_300 : v3_1489577445_306;
   assign v3_1489577445_306 = v3_1489577445_307;
   assign v3_1489577445_307 = v3_1489577445_19 - v3_1489577445_46;
   assign v3_1489577445_308 = v3_1489577445_58 ? v3_1489577445_309 : v3_1489577445_300;
   assign v3_1489577445_309 = v3_1489577445_315 ? v3_1489577445_314 : v3_1489577445_310;
   assign v3_1489577445_310 = v3_1489577445_313;
   assign v3_1489577445_311 = v3_1489577445_312;
   assign v3_1489577445_312 = {v3_1489577445_217, coinInNTD_50};
   assign v3_1489577445_313 = v3_1489577445_19 + v3_1489577445_311;
   assign v3_1489577445_314 = 3'b111; 
   assign v3_1489577445_315 = v3_1489577445_316 >= v3_1489577445_322;
   assign v3_1489577445_316 = v3_1489577445_321;
   assign v3_1489577445_317 = v3_1489577445_318;
   assign v3_1489577445_318 = {v3_1489577445_217, v3_1489577445_19};
   assign v3_1489577445_319 = v3_1489577445_320;
   assign v3_1489577445_320 = {v3_1489577445_52, coinInNTD_50};
   assign v3_1489577445_321 = v3_1489577445_317 + v3_1489577445_319;
   assign v3_1489577445_322 = 4'b0111; 
   assign v3_1489577445_323 = v3_1489577445_324;
   assign v3_1489577445_324 = 3'b010; 
   assign v3_1489577445_325 = 3'b000; 
   assign v3_1489577445_326 = v3_1489577445_62 ? v3_1489577445_356 : v3_1489577445_327;
   assign v3_1489577445_327 = v3_1489577445_328;
   assign v3_1489577445_328 = v3_1489577445_60 ? v3_1489577445_343 : v3_1489577445_329;
   assign v3_1489577445_329 = v3_1489577445_55 ? v3_1489577445_335 : v3_1489577445_330;
   assign v3_1489577445_330 = v3_1489577445_53 ? v3_1489577445_335 : v3_1489577445_331;
   assign v3_1489577445_331 = v3_1489577445_51 ? v3_1489577445_335 : v3_1489577445_332;
   assign v3_1489577445_332 = v3_1489577445_41 ? v3_1489577445_339 : v3_1489577445_333;
   assign v3_1489577445_333 = v3_1489577445_39 ? v3_1489577445_335 : v3_1489577445_334;
   assign v3_1489577445_334 = v3_1489577445_37 ? v3_1489577445_336 : v3_1489577445_335;
   assign v3_1489577445_335 = v3_1489577445_20;
   assign v3_1489577445_336 = v3_1489577445_36 ? v3_1489577445_337 : v3_1489577445_335;
   assign v3_1489577445_337 = v3_1489577445_338;
   assign v3_1489577445_338 = v3_1489577445_20 + v3_1489577445_9;
   assign v3_1489577445_339 = v3_1489577445_81 ? v3_1489577445_340 : v3_1489577445_335;
   assign v3_1489577445_340 = v3_1489577445_80 ? v3_1489577445_335 : v3_1489577445_341;
   assign v3_1489577445_341 = v3_1489577445_342;
   assign v3_1489577445_342 = v3_1489577445_20 - v3_1489577445_46;
   assign v3_1489577445_343 = v3_1489577445_58 ? v3_1489577445_344 : v3_1489577445_335;
   assign v3_1489577445_344 = v3_1489577445_349 ? v3_1489577445_314 : v3_1489577445_345;
   assign v3_1489577445_345 = v3_1489577445_348;
   assign v3_1489577445_346 = v3_1489577445_347;
   assign v3_1489577445_347 = {v3_1489577445_217, coinInNTD_10};
   assign v3_1489577445_348 = v3_1489577445_20 + v3_1489577445_346;
   assign v3_1489577445_349 = v3_1489577445_350 >= v3_1489577445_322;
   assign v3_1489577445_350 = v3_1489577445_355;
   assign v3_1489577445_351 = v3_1489577445_352;
   assign v3_1489577445_352 = {v3_1489577445_217, v3_1489577445_20};
   assign v3_1489577445_353 = v3_1489577445_354;
   assign v3_1489577445_354 = {v3_1489577445_52, coinInNTD_10};
   assign v3_1489577445_355 = v3_1489577445_351 + v3_1489577445_353;
   assign v3_1489577445_356 = v3_1489577445_324;
   assign v3_1489577445_357 = 3'b000; 
   assign v3_1489577445_358 = v3_1489577445_62 ? v3_1489577445_386 : v3_1489577445_359;
   assign v3_1489577445_359 = v3_1489577445_360;
   assign v3_1489577445_360 = v3_1489577445_60 ? v3_1489577445_373 : v3_1489577445_361;
   assign v3_1489577445_361 = v3_1489577445_55 ? v3_1489577445_367 : v3_1489577445_362;
   assign v3_1489577445_362 = v3_1489577445_53 ? v3_1489577445_367 : v3_1489577445_363;
   assign v3_1489577445_363 = v3_1489577445_51 ? v3_1489577445_367 : v3_1489577445_364;
   assign v3_1489577445_364 = v3_1489577445_41 ? v3_1489577445_367 : v3_1489577445_365;
   assign v3_1489577445_365 = v3_1489577445_39 ? v3_1489577445_367 : v3_1489577445_366;
   assign v3_1489577445_366 = v3_1489577445_37 ? v3_1489577445_368 : v3_1489577445_367;
   assign v3_1489577445_367 = v3_1489577445_21;
   assign v3_1489577445_368 = v3_1489577445_36 ? v3_1489577445_371 : v3_1489577445_369;
   assign v3_1489577445_369 = v3_1489577445_370;
   assign v3_1489577445_370 = v3_1489577445_21 - v3_1489577445_46;
   assign v3_1489577445_371 = v3_1489577445_372;
   assign v3_1489577445_372 = v3_1489577445_21 + v3_1489577445_11;
   assign v3_1489577445_373 = v3_1489577445_58 ? v3_1489577445_374 : v3_1489577445_367;
   assign v3_1489577445_374 = v3_1489577445_379 ? v3_1489577445_314 : v3_1489577445_375;
   assign v3_1489577445_375 = v3_1489577445_378;
   assign v3_1489577445_376 = v3_1489577445_377;
   assign v3_1489577445_377 = {v3_1489577445_217, coinInNTD_1};
   assign v3_1489577445_378 = v3_1489577445_21 + v3_1489577445_376;
   assign v3_1489577445_379 = v3_1489577445_380 >= v3_1489577445_322;
   assign v3_1489577445_380 = v3_1489577445_385;
   assign v3_1489577445_381 = v3_1489577445_382;
   assign v3_1489577445_382 = {v3_1489577445_217, v3_1489577445_21};
   assign v3_1489577445_383 = v3_1489577445_384;
   assign v3_1489577445_384 = {v3_1489577445_52, coinInNTD_1};
   assign v3_1489577445_385 = v3_1489577445_381 + v3_1489577445_383;
   assign v3_1489577445_386 = v3_1489577445_324;
   assign v3_1489577445_387 = 3'b000; 
   assign v3_1489577445_388 = v3_1489577445_62 ? v3_1489577445_418 : v3_1489577445_389;
   assign v3_1489577445_389 = v3_1489577445_390;
   assign v3_1489577445_390 = v3_1489577445_60 ? v3_1489577445_405 : v3_1489577445_391;
   assign v3_1489577445_391 = v3_1489577445_55 ? v3_1489577445_397 : v3_1489577445_392;
   assign v3_1489577445_392 = v3_1489577445_53 ? v3_1489577445_397 : v3_1489577445_393;
   assign v3_1489577445_393 = v3_1489577445_51 ? v3_1489577445_397 : v3_1489577445_394;
   assign v3_1489577445_394 = v3_1489577445_41 ? v3_1489577445_397 : v3_1489577445_395;
   assign v3_1489577445_395 = v3_1489577445_39 ? v3_1489577445_401 : v3_1489577445_396;
   assign v3_1489577445_396 = v3_1489577445_37 ? v3_1489577445_398 : v3_1489577445_397;
   assign v3_1489577445_397 = v3_1489577445_22;
   assign v3_1489577445_398 = v3_1489577445_36 ? v3_1489577445_399 : v3_1489577445_397;
   assign v3_1489577445_399 = v3_1489577445_400;
   assign v3_1489577445_400 = v3_1489577445_22 + v3_1489577445_10;
   assign v3_1489577445_401 = v3_1489577445_105 ? v3_1489577445_402 : v3_1489577445_397;
   assign v3_1489577445_402 = v3_1489577445_104 ? v3_1489577445_397 : v3_1489577445_403;
   assign v3_1489577445_403 = v3_1489577445_404;
   assign v3_1489577445_404 = v3_1489577445_22 - v3_1489577445_46;
   assign v3_1489577445_405 = v3_1489577445_58 ? v3_1489577445_406 : v3_1489577445_397;
   assign v3_1489577445_406 = v3_1489577445_411 ? v3_1489577445_314 : v3_1489577445_407;
   assign v3_1489577445_407 = v3_1489577445_410;
   assign v3_1489577445_408 = v3_1489577445_409;
   assign v3_1489577445_409 = {v3_1489577445_217, coinInNTD_5};
   assign v3_1489577445_410 = v3_1489577445_22 + v3_1489577445_408;
   assign v3_1489577445_411 = v3_1489577445_412 >= v3_1489577445_322;
   assign v3_1489577445_412 = v3_1489577445_417;
   assign v3_1489577445_413 = v3_1489577445_414;
   assign v3_1489577445_414 = {v3_1489577445_217, v3_1489577445_22};
   assign v3_1489577445_415 = v3_1489577445_416;
   assign v3_1489577445_416 = {v3_1489577445_52, coinInNTD_5};
   assign v3_1489577445_417 = v3_1489577445_413 + v3_1489577445_415;
   assign v3_1489577445_418 = v3_1489577445_324;
   assign v3_1489577445_419 = 3'b000; 
   assign v3_1489577445_420 = v3_1489577445_451;
   assign v3_1489577445_421 = v3_1489577445_425;
   assign v3_1489577445_422 = v3_1489577445_423;
   assign v3_1489577445_423 = v3_1489577445_14 & v3_1489577445_55;
   assign v3_1489577445_424 = v3_1489577445_12 == v3_1489577445_52;
   assign v3_1489577445_425 = v3_1489577445_422 & v3_1489577445_424;
   assign v3_1489577445_426 = ~v3_1489577445_427;
   assign v3_1489577445_427 = v3_1489577445_428 == v3_1489577445_15;
   assign v3_1489577445_428 = v3_1489577445_450;
   assign v3_1489577445_429 = v3_1489577445_445;
   assign v3_1489577445_430 = v3_1489577445_440;
   assign v3_1489577445_431 = v3_1489577445_435;
   assign v3_1489577445_432 = v3_1489577445_434;
   assign v3_1489577445_433 = 5'b00000; 
   assign v3_1489577445_434 = {v3_1489577445_433, v3_1489577445_8};
   assign v3_1489577445_435 = v3_1489577445_50 * v3_1489577445_432;
   assign v3_1489577445_436 = v3_1489577445_439;
   assign v3_1489577445_437 = v3_1489577445_438;
   assign v3_1489577445_438 = {v3_1489577445_433, v3_1489577445_9};
   assign v3_1489577445_439 = v3_1489577445_82 * v3_1489577445_437;
   assign v3_1489577445_440 = v3_1489577445_431 + v3_1489577445_436;
   assign v3_1489577445_441 = v3_1489577445_444;
   assign v3_1489577445_442 = v3_1489577445_443;
   assign v3_1489577445_443 = {v3_1489577445_433, v3_1489577445_10};
   assign v3_1489577445_444 = v3_1489577445_106 * v3_1489577445_442;
   assign v3_1489577445_445 = v3_1489577445_430 + v3_1489577445_441;
   assign v3_1489577445_446 = v3_1489577445_449;
   assign v3_1489577445_447 = v3_1489577445_448;
   assign v3_1489577445_448 = {v3_1489577445_433, v3_1489577445_11};
   assign v3_1489577445_449 = v3_1489577445_38 * v3_1489577445_447;
   assign v3_1489577445_450 = v3_1489577445_429 + v3_1489577445_446;
   assign v3_1489577445_451 = v3_1489577445_421 & v3_1489577445_426;

   // Output Net Assignments
   assign p = v3_1489577445_420;
   assign coinOutNTD_50 = v3_1489577445_8;
   assign coinOutNTD_10 = v3_1489577445_9;
   assign coinOutNTD_5 = v3_1489577445_10;
   assign coinOutNTD_1 = v3_1489577445_11;
   assign itemTypeOut = v3_1489577445_12;
   assign serviceTypeOut = v3_1489577445_13;

   // Non-blocking Assignments
   always @ (posedge clk) begin
      v3_1489577445_8 <= v3_1489577445_23;
      v3_1489577445_9 <= v3_1489577445_64;
      v3_1489577445_10 <= v3_1489577445_88;
      v3_1489577445_11 <= v3_1489577445_112;
      v3_1489577445_12 <= v3_1489577445_131;
      v3_1489577445_13 <= v3_1489577445_152;
      v3_1489577445_14 <= v3_1489577445_170;
      v3_1489577445_15 <= v3_1489577445_175;
      v3_1489577445_16 <= v3_1489577445_206;
      v3_1489577445_17 <= v3_1489577445_220;
      v3_1489577445_18 <= v3_1489577445_249;
      v3_1489577445_19 <= v3_1489577445_291;
      v3_1489577445_20 <= v3_1489577445_326;
      v3_1489577445_21 <= v3_1489577445_358;
      v3_1489577445_22 <= v3_1489577445_388;
   end
endmodule
